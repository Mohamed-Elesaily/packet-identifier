module decoder_64(
    input   [511:0]data_in,
    input   [63:0]DK,
    output  [191:0]type
);


always @* 
begin
    
end
    
endmodule